[aimspice]
[description]
1783
testbench

.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 3m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R2 NRE_R2 0 dc 0  pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

X11 1 0 EXPOSE ERASE NRE_R1 OUT1 OUT_SAMPLED1 pixelcircuit
X12 1 0 EXPOSE ERASE NRE_R1 OUT2 N12 pixelcircuit
X21 1 0 EXPOSE ERASE NRE_R2 OUT1 N21 pixelcircuit
X22 1 0 EXPOSE ERASE NRE_R2 OUT2 N22 pixelcircuit
Xmc1 1 0 OUT1 activeLoad
Xmc2 1 0 OUT2 activeLoad

.plot V(OUT1) V(OUT2) ! signals going to ADC
.plot V(EXPOSE) V(NRE_R1) V(NRE_R2) V(ERASE)
.plot V(OUT_SAMPLED1)

.include C:\Users\Jonas\Documents\Uni\19W\design_of_integrated_circuits\project\PixelCircuit.txt
.include C:\Users\Jonas\Documents\Uni\19W\design_of_integrated_circuits\project\p18_cmos_models.inc
.include C:\Users\Jonas\Documents\Uni\19W\design_of_integrated_circuits\project\p18_model_card.inc

[tran]
1n
60m
X
X
0
[ana]
4 0
[end]
